module ADDER_4 (

//input data
input [7:0] PC,
input [2:0] CONST,

//output signal
output reg [7:0] out_adder);

CONST = 3'h4 //adiciona 4 ao indereco levando para a proxima instrucao
always@(*)
	out_adder = 
	
endmodule
